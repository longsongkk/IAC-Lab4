module task3 #(
    input logic []
)